Circuito do trabalho prático
V Fonte_1 1 0 24
V Fonte_2 3 0 15
R Resistencia_1 1 2 10000
R Resistencia_2 2 3 8100
R Resistencia_3 2 0 4700
.END